
package yapp_pkg;

    // import UVM and include UVM macros
    import uvm_pkg::*;
    `include "uvm_macros.svh" 

    // include my yapp_packet into package
    `include "yapp_packet.sv"

endpackage : yapp_pkg
