
package yapp_pkg;

  // import UVM and include UVM macros
  import uvm_pkg::*;
  `include "uvm_macros.svh" 
  // include my yapp_packet into package
  
  `include "yapp_packet.sv"
  `include "yapp_tx_monitor.sv"
  `include "yapp_tx_sequencer.sv"
  `include "yapp_tx_seqs.sv"
  `include "yapp_tx_driver.sv"
  `include "yapp_tx_agent.sv"
  `include "yapp_env.sv"
endpackage : yapp_pkg
